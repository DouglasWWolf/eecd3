
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
//     This module is used to narrow the width of an AXI stream in order to trim-off unused bits
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~

//===================================================================================================
//                            ------->  Revision History  <------
//===================================================================================================
//
//   Date     Who   Ver  Changes
//===================================================================================================
// 14-Feb-22  DWW  1000  Initial creation
//===================================================================================================


module axis512_to_256
(
    input clk,

    //========================  AXI Stream interface for the input side  ============================
    input[511:0]    AXIS_RX_TDATA,
    input           AXIS_RX_TVALID,
    output          AXIS_RX_TREADY,
    //===============================================================================================


    //========================  AXI Stream interface for the output side  ===========================
    output[255:0]  AXIS_TX_TDATA,
    output         AXIS_TX_TVALID,
    input          AXIS_TX_TREADY
    //===============================================================================================

);

assign  AXIS_TX_TDATA[255:0]  = AXIS_RX_TDATA[255:0];
assign  AXIS_TX_TVALID        = AXIS_RX_TVALID;
assign  AXIS_RX_TREADY        = AXIS_TX_TREADY;

endmodule